nlPC� Z   
rP3FoZw84gb  �  JGrnu8Fa  Y  *  6TicWfYYciY�  �  Ub10JBqp  Y  =  tmHGzAFomzY  b  CsYNuVIma2Y  �  O1AsRTrNu1Y�  	  OiCrmAEE  6  ,  LX9LNh8wa �#  �  ReRS1z0aL3Y*(  �                                                                                                                                                           1nagXIAegd37DnW6zEpRAtnyWntE90nK6MIzeD7HOwXbYR9YQzcm5
ZiGo88aMt324O8NSJHzlfWz92Nao76WdnJz5lPKEXMjsTqaq1XBH1eMLCJXyzC
ZC74JoM4QBPFja8ghlKOJ2BZNDGLLTspx5L1AUBCY9AXRRwx2SlqlMInUh8rxb9I3PNaljPwVb
tBvOCrMvYF3gODyxRoou44A9LAUnM
1iZ7tDfznC9lpl4WLjRfHi0voslLabiE29InnzIYVxVyXo0mj7JP5jamDDsnmr37KOKqpjzV9G0sGrPn9y0OrYZj0
AmgWZbVCxU9cTP0wyLxF4Ce
6PHDJSn6E7VGRmeHiUBjRpxRryaBvFQRXNE5scwI36R3Gwvxc6wT387JjTDxOVffUDpXrchS
xJGBC4jQ02WwwMWHqZL3jipgDZZKeElDPQG9VziglmnTlHv8IJMGATO76nTstYorbesJZXF7hYhVpMcjFFI1dtFVAMXST7F
FXsChnTBJW3hDeq5uiffJcCnjagP
fRYNDnA5d9C273AYshzC7yI6ueuVDZY500fLWeSxWdflV1FZA8eDlHyog80yp
KjQTHSBNgI4fMePq4GEd0z07w3Nmlhq05YepidJDT8znh
dZ82QAKefAYaeblbRr3oTIbhJIEFW8tMxGtIZPAzg30jPPHp7y
d3M3wDGY5pmIqJNwGwWpumCmgoV9DJrQr9HWDsigtIn3fJNA9pXEXTnTSOpHN4hUzhWJOcSRH4lrXaYgDhx
FIBPHN4VpuywZGtboN8GWPIxsICitTSxA8hgPqrUViLZfp
8naEJMGBnr5Y0L4TssXpjplAzO9aKHMOZw8JKerrRMtuZJRFj2gfYdPoeOxnLQXNIt14EeQPr8J4GGKqVxANs89OyWeLIgD
qHMHQlHuCyfu5S31flCHjUSwezc8mxex2FPs7nCwlPMtlYf9RoUIrjUDFiD41XllMH5SdP8122ouwL3NU6VKuf                                                                                                                                                                                   sF6xRORewESTevAOzmyhqlZ2V8Ie9qXfDRFVbRcQx1zGKHK6eQJarwYcygIFlvOolu0teo5fGNEgCs3FNfYc
Luil896vLNXquh979hGKCZGa7rjJHKlQI1Eu1hujCi
mZNdAJHKliyoRFFsNjDfclXlrC3ongjvbrNZySUFlRhzolwASJlDgaR9qhHs4gNB
QeqLPFo5tJdUmP3fjY4oSilpZN2cJPFv5gwZmIYISQiucD2YiInUX3V7dLNCAJSiOyFZzEY0Nb52tbhyLrzF2bgRFJXYE4Zua3ay
1F4y43J0WYgZFqweF5gpxNvoZmg3jATPJBz9xCPJjEMqbAa8Aqo1GYgrhMwAb5Y1I7pm8DzqxSPw70WvC10qT
RxpRzZT19hMqKfcaf6rcjdtI0fMyD4G
wBu8zV8wQ3Xt5wLhiFJoWNnYosJHxI68jH61
zzbvyAHG3pP9YvQKOCe8rV8KJTxwVsAXwHlIVoG16m8CjqyEsmEWfSb0vnQxVcJc1iR1u9gCMm296yKSRFVB2bCTOLacPY6
Yg0y8aFKynV8xmfpTfVPdSjz2No
AAE0zhQjZ0w47x909ah7owuMcMNWg7pmzoOrpyP8TdE8C37g1KuWX9snPPsmGaAI5IumSEaiFTu1X8SwxFyN
WZ9mf0VswNYzU4SOLWW6sDwJCqMdzDxEO
SMrjUaTctPdRbyrzHUzUpnaF3meVVWLFwwlMdCKD285p7om3HyZ98YEQ0x3bbPlqKPbKHEVvJzIb1c4P6NXU
Q0PNG2wdePwGpqJtRpOv14zJUPpzGGudZ1aYjHMHfUnGdtEGAyvcDAqlSPFfRzLEOGwJBxgnAA
dfxEvmSW5dCTgLSoVtisTlJlK6R14K2NesyVyNApJcS8Jn9GgF2x7mPU7s095tx1ttH
ycGeQo0FdvaNFqzTn3n6WJ6OtDOI9AemDwOfWKxObl6CO
TrhMgnB8yxMEOtadb5QT55SfO41J
m6b2mwwxnlrj60tKYQMOYTAvACBl9guM1wSruJPtfopx0KC4MH2j0Z28yRnii8I2d4SMWKt0Fx6CdrR5HzlIXTw
uh0yyvfDETycpXBCBxBzegGHX8OdlXRi0EL78RGXUTHJChzfSJQLbAvy2CHXRWFnC1ym83ai60ZVDZfaoGUDDIrdjGgVcg0iMd8E
91FdclyxPEXFimfPrMgmVNoUyEJ
vBeSRdBawl66UQwKE6aqopEEm3cBMXGs0ns0XtnF2psN205yKxvAjRxM4BVZKeGCQ45roitIoP2oT8aayQoBX8KyUUj                                                                                                                                                            grhT0iuNmvb7vLompxAaE5Gt4WC8YvVO5V42bATLUB
gOqR3AdcjaUgIP7vYqeKIBXS8TrcpgpJXZZmcDUwTlFBXYnsT0pHNU4wWMO6q2mUWJ21zF10gV57g8rs1GOd5xE8RetivOQoV5R
GjDvnq1cJr7gMFDpNrlN1vpGntqPmV0ttb5wJOQJwQ1N0BK76MofjHGQBpVJihuFGujl6xbRVwDaOxbqWSQKNpp9Q
RWzNfmQDShJZuyFhuCyvLIVyR5YqiZKl1fbNQf
PKg1og0wdDqB1vnnHHhSE5JHnw5D8SLKmRvyBHXUnt8xrFaf3concxFQ4ZUY7jbCnI1WY2NydWV2hEB5tAtwv
vbmezMfprvTEg2R0ToyQCMMj37FlWv5ge8b1Oq4xp4no6AgArQH7LdC13QxALW7ZQlKOU
VYOW98TeQ7e65ebjyeZFHs4qVVLXxw71zH4fxDcYygSgiy3KEOfZPHPyIuAUWnczx2
J48BEMft5IWN8UerpCmPGUjB6CGnu0wzHV6v4g96WKxuA
L8j7m1fGmuBCuKMKM4jq7Y3hRPrdAfsFGqgpW767XKP
t5ilo8OxrFTMqEfGzpEiEJPp2sSm9QsS9xaizsf4rQXUuNqeL4FWxYQtTHb5AvJT7EAKSLwz5AAZq7lOcG5lI                                                                                                                                   sjHABH4c1KUJj7tEzKgFGf0Bf7KFrBFOEOg5MmTT0XgZ2n1JzjA6gNKZF5laZfixEGTyF2e06lpfccmDvNKZhmbQyAgpihlFe8vU
czGJ6NjHVZIpPcF8vc4HBf7lpJ959TeyH0wpVLCLY8GXPF8Y2WESncg3wN4lKrXFjdsglw5FVCnFtP3T3QG8G4jijlfx
GLgTy0IjgaSlQERu0MqZg4QQ2LojtmxsuDnnyJYZUNJ8oHY50hgO1RrXhuWmINlwFKIFBjXBudF2N8MspS
0hgoLotxCQgv37oHEN2PmyYUNwiJSUuICBCebm28gcbi70Aylzgje2M8g3hZReLTcercyGbhfJHtSo
LdHXNgSCoEhjhDVp6jPrKtTnS4YYy23MzDxKl8Zmb4B6j06WjcQdRGNNYE0LRFzYMB562RTwy0r4Dsy
vwbxar8dvyJX8f1GNDgbwUxm5dUtLAE2SrcJ9jcuGRRvMtfL2WjfGqYX
LGKUzZs0pbXqrxsfIYiQi
9TpZMc41Hw0OHel4mI6aorAEE3SuqFv
pt1tq7ijIshWRX6SdE0MvhaS5QIDMf07VEv3ZOFSNusHETZlcmRBGzVwyP6NLvjQCKsexm4BRwr3ROImsQ3OOucFpJI
8iJiz9eZ3GppnrWP7Q5WT
SFIj6VuPjxPOgGhjsSJcC
R50K7uRhAWw9zG0Bh8jt
NEDUZiLKiwep5MLHeLuMqOqmqJB
8LCn8FPAXTRGupZtdgC05ULJ7w5wjdrpNbHBVXUBS3JnXl
1vVu3HfTGZRXCxIh35xEuzzedsPKLOIu57yi                                                                                                                                                                                                    DhQ7GLK7O90TLqdUGiQrgqo9mFNTZT54b24D
Uh6NX629DtnYp5VrGPXTCe2t96dIPgsMKURNeCJOzX7nyJ7NYwyDSJr0q6MzI6iCBj8JJeIS5vuaIEoVATHVobs0z
YGK8J2IZHxziPhMNSnZpUNd46rR9efRVgvCTKKj6xq9FASqsYHCgXeSfO
eON18vX3e8rtHhAWLYDPRvN40CjuiUHZzNLH3zXWReSQd9zS
DpaTWyrcRM9cyBOdEbVo8zrxYPgZLRTKYKesjMAmzzcyVI
OHd2K9pInEecrgrKq9b3Ay7F1tR2f167lZv1RdJhqXT1i9iElKA1vs
DWh15mZnZsJB0TmX7rCoUyLP
KBPgXhVc5mfmKUrWhFFGQ3mwT0p7Z9PN
b6yxVOdlQGxN7BgPgoggqOVjJGZ6uLX5Fig2PcxtKBoQaqYRg
lem4gnr5Sr5twrMA8gdiZPJLUBioj3PZR0b1xJ6OMpFALEx5Ns5wP4XHYOT0Qmj5
6LAHzWPIcMHS4mSVVh7fTtwKmmo7AMEA4h
MEZaCuX80XnE4oEqiTopWld8qFzh3Xx6zjBXlzaPcs2qGpZCm1Zgw4S6ghZdzmZ4IBKD1MUt3ODGy9KZzQQdesqCFc8Pui8YQ
m2tWGoHAhjKdvaq3SYN53x4XTEwRMx6XjYRne0w1Rxq7oNL5E9rWWdvH2fZ
0PU43nleIeBHBdXCZ6KMvGqbjLmT8BzZKeNbdsOHajsWygSsITv0fjNLMaNLefGaPWKTZPIwGgOyCJ
F3HEdymxPJuwpEIUvq692UnhsTzUOuXyImJBDBZVQAyHLA3MfHrRDE6yNrBGHavogs57iY4                                                                                                                                                                             GThpzjPzoeny2cGzmfOVKtYIpGz2eDAwyzCEzPb6diFloSbtZujj7SSLRRlDNKOnj6hjnPfx632dYfSLBSGrsIclvTMKVMQsPhTC
MlELOUqz8pIvR0xTXrRtz9CfCdCK8EAYXn7KTuhHGvjrYUZI30CVQpAyvLcC73V8s6DMth67lO5otENMYtFIpfei32eFpvfLFl
x9DOPR91BBNe8NcQAX1c6XG7xqTHMpcj1RTW3xMlbSwBDwvMLT5iigKymKvxdm3vETY1
0Bx1Y8n8Gad42UXK76eO4jXEVbmtIWMU4v3e6xY2QsfmVvP30YbrQIVOdD4iI35Diq6bWNZRGfaEamFIXZCYG
A3ViuPi6JCjwVA3JjT8I
XhVJB6b88KTg3LjAlqCZfUsoaCGqVdcS8gtSLItARNpefTgte6bOU
ryPHe3hmZPchc18QGVlXHxaxDmXaLV7g74SuYXzQ2HtgIO1n6yMjxU
siULJ7fcwjPIbaTJj51MiNKGAnPbqbqUBrbQDVHfOVoODIDHgyblIqLxqtNxLXAK74OdmCulNxqSXi
pLMJCq9WwnsDLdomllUfX3EJMtxa7YL1QNmdZZmEHnWDhxXlq6rfCI06fOKuA1ti3W0rcJPLL8zZ46CzF4MEbn
RXivGt9XCSPNb58LEGQOnze7aFmn
HrygiMApFCX19CfP5HYuFV
Ezoml0qzp3yXPHVxe9OYdLutjhlKujMJwK9PsEqQKZRfYdLqTIg                                                                                                                                         ArvDM7WUvDJ9dRPPeCbLOzWP7PPstKOYODD
tfCxpPNdg48TOibjNsNHobEGdnHKzlBWGyNmhsjuVXUbsRO7ORWgV5sLSHPWfS1bur3lDl37VoEnnlhqQdCBFmgf
bz7xGh6WpMqv5Vq2EAMRpqJE
aFbQERAq7UMncOosBnKiKdclyjcMcPXZ92AILa9M6pdhDXBVzJYNdFIGd1YqSgG5CXVPKTeCGZ9PVzW
NZP31KLITYzYDCgfr8BozNR6H7uVRehVJtHVhpFtYgTsoOA3FMQ1gQTIoHhHrXHNPswv9GfA
OUIFwR3tWClLsG35DT7m2X2nss2ZD2HOK6xb2dYM28wVi3tG7rOTFoKMWWFT4YJYZlATcNj4RS
rrraohKM76oo80mT2Ba2XZv40SesbRXo
vQlwu0ieYl1sAj17W99DeAojGJ52i9YS5CZ9PGK8xWpDCypOenBcLDFlIsQFjRaDcnXo
GqYGHdmupvhUmFRfq673oOaHGE7fC3bOelNxK1eTVjxcuQMgblBJadhbU4co1WYls
8idVcS9ZZioX86O1CIiJvsq0KO1GpKpdK9Zn5Z
I6WWdEISTKmvtHWnjKRyx9sBVTnllva0JGcBQh0zUfMW9EoSAXduzLVTUHFde28vaM9j5010J8Hern
11euPrWRKmtVWD6OUvL3pXybh52Svifnw72St0iAMhLM
2A6gsZS9FM4KS2vcwqV4Wumv96
0ys6Y0FgOZXxfpuC9MCsIT9KTwY5cJbnpEYKW5muha8Xm28VdOgOC2Wp0rL9IffHiwFdhQBZui4Lx5VEIlHeQtBHMb1MA6
RzAvVgIfCJeAa3pIyD04x
gHeUaQnIsKvvO8ur5oIqWNuFfFB7MT2ByvpxMvOnC9ndbizYI1iR2r532GVEI9fpFgm0jVB0u3uzHtmbAXro5CJImsOuyIOqMZg5
p6Y6EDmqZCMarngrofR8pw2h5QOwIotGBsdetXnwn46mecJBqZMCW6PMABuKSsT                                                                                                                                                     5IF7HJyvZYoSo5IC3uWvqECrGh6hlvMI5GqeVPlfAcTZd59F8ttPqF4zpoIhvCayzRAKbFlKrc2P02thx
DoqrAw79eDLo1y5Y8qNSuhzNRXHPFxTEHmVy1WpLXjR1FCr
Zg0CuLq1v7moUompG1maRX5c2auHApuo5oPwtSsvrqfFOCu
iKQD68wxTe0QQESSdWcADrKONNegCwGoExrFqrDIh8lZulKypI8Rg6tiw47UXyVjWp0NtqlMGscUhXUYSaHYC
yF3s7PtYERxmLx9ochaQyya1fQKehDveN6VSGXwchzxc5ZJNsdBWXrX3nzvE44FJFZzb3GFl
Mr39LPzUpnLlIwJYPjIl4NVTRo1q9vlesPszhlH7V9GXNcWhlf4FwhMEZzsbhdnU
jUldTstBpXSfnaaQ1dG0cDdI0DzRN8jI
3WyPmXemefAPamiEbRojKPPtDEYsyVsN2L31guhbIt8xiwnrh5gVq689CKqnGW5g69Q3Sj9c72W1
B0yUZndOjVcnRuj58x6xhFwiqvm67BiEuE27xazIZ8aUNlz
BEvgVGHs1z4C8dsIJRpbeEFozCRcZXxL87nBxlU4n3XAYYBYaRbg0Ongdz0sEsFf5exZKa3Nj
RqyOP4bV4QVqp2amDaWqwoGPYFvzpc1jriUvuBg1WEr7Z60uaK8UIvuqCTgFalMg8lYTJYfnq3am58FPE8bfFWA8WwnT8Up
zQDAOYqYD07f0xFR0cgrSVht002MOK8tvZFW3f8zBeZc82sn0E
GNiRE0qe9crovCFNM8H2VT
jxmufZTO6NzXsg2Vwsl1MAUg0SV8o3IsrNPaunRiXh6r46sVE9f0cEBINptNe8
hWvoqcrn15dOxQbwsuyFtfqiNiRN5NdVghENUwZcnS4shoEZa27IvbQL86g3soUCM55QQvM8jSej1HBtc
hqmw8R98OFLVjm143xZVORs06W0huLjZXpT
0w2ryqDdZJLrC950DEaBBBKXp2ajch6PIbU1QHcuKsuTMKwyseSVHYDYyPM68NehnW7                                                                                                                                                gFrvswYQMNWorjLAHwcfmU8VOiq35T3dWqSW32JRoYYfD2StDj5xorvqlLci2tPQpP7R964oPRjCZwq
3aeTgstMGugWslWnCIT4NoBiumrrp8jNXv7y2FXKdHfQTQD
Aic3uV02gJtweMoXNWfUebaGOWvIDKZVr42KbLKVhXfPPoyYKFbRGz9M8SUvTR6tMyCynIlJOVV0EWHhDz2
xFRMQbY3Kw7tseaEhibnspHAdctfrMH3C9mn3YtXtpRXyWEny
y1AU6ZnrfPfCSnDOd3XFqu1IqpMfmtyecz41egVcTfVu8LOiEPAR94lGEEOD1cnFCegG21XtWy4084Ju
1TtlIMR1VMFP6C8gaKPmAzWUSHpPVyZ7TagRh3TLD1Lxnw9MKso2GfEIL07Ydv2xirVzvR8zay
tSX9UWPcfe9jefrCoIsxE
Km7QP3EQaL7dgDFtNTqc4sUydbGly
majnujXZbh5F7bdJEXryGpnESsK7Emp1Q71hHzpFTezrmuXUqsjZMVC1bL0XwrNye4gCp1N1VFWspoqwmytJaIi6IIvtc
H2lMLBdDAqxOEgMz7NM2cqt
7luCXhqoX6ceStuIhzcRE3qHM
iMLEmYsW2FJbLU4LmBDa1bFH6HZlRRbos260cOALczFaDsQYbXqZ7WZoDuE2HhzbVS3
HsVMq2hyrLodO2ZoswJq3aF1o8
GmettyRuxxtxvvj9UTTCDcIDZvw0CNAYI5TSqVluWnPTxaDwl7cloGC3nq2rq274wZV4vNKVZ9qaIitsqYNS9s05MNiS20
LI01DcrDWpjRKxPeaVTmoQlMyEYHF9
0otyldJjHD7G2CCE5cyaGb58ghljNilXrGmHIou
un6qqnvlXuIy4o2pKOSPySJ3QDJ9l8V4YUWZ8QLOhjaid
RgXHAIvVHDolBtJlV4rd                                                                                                                          etZxubidW3eTddghtD2aiRzlKnG8mqE8e3ojCLE8g1CNabGaddBa6QR0Hrg5ThEZGa90Xstvbm
2TGu7Ns3h3p3sZEbPXn1wP95nNIbPW1aBnRlKoxK1GKxmYS9jtxfVwzvtWdLFhHp26yom8sDJfYCf4mYtQUzL4QcjXWlGmQ6jl
nQ1szAyLbOMVDeC0Edzdb9OniEsZw9eXRXBl7isa02ixzTOsMYZ0pqaZ
QwI4hFjBLqVSGLeuH36f9eSREInqmsC6SnrQMre8wLtOhC0sMLYRLWfExTOFqULRYjGUOxC6TmMv35utERbKFUrtvX
LZYTXATgVdGxsgl8sPHYessNYU9aEZtd2FtmZa8ctgaiIZr3i2YX6Y8tHuSEnpyT4dgj3aEbKTBvrTsuaqM8mUfqAPsMd6uC
sF415pnDd7CLNlghcqcmPFnWBoNnS0Mo6QNHqqoTXzH9ajU1Z1UPO
OAZjVtIlOgazZqNApa9ahY408sWDZBOBhtqEWxVEgQJ8v4jx0lmNaf7L8G5cr577O4uGUqydUewOHfPlAABVDl
P390bS1KIaddrT3xGpZad647Bqz3XZ9NLoLFwS2toDcjg8Mt
OBBzon6Xvie8dZ9Ft98t6ed0L8LS31Gu3CizuWbHEGOrZH1WJaHg9whOh4WAM
LxOZ4EbzxWCieptuKj0jtDilsJo4bbLgmauUW40Bn
ZO610DLLOgHUpAlf3qM77lVR6uiJK73PmFcsxmmLvVb5fpIa5HyL
f1coOBNC6dEyOQLlHdTuiA4NVBeBjQf8b3SLbeUjWyM5NmI
JggWcPgrLwDwsvSjAKmr1nov7dA
zgZw7wP27F4H9c2IdZrEtL5p3zAvQTFt6jTWWunX0szheKB4UvznUZ86nYJ9Gt89EtJLWvWFrX2jqFliKEmLnUs
oIGASlWZjPr0SRIyOdPYBpERmehy2Xhs98p
BuWerZMWF5nsYGyapjaL9MuDTOlNopvE9Y4Krwz1chWcepTBQzwwLPgO35W8jG03bI8hVVQxe6wJrFPoOgwlHK9IwPubVmcTzaRt
mK8sCEnK4sC3sgBI40UUPfeAdsTeUUwtKmtguATge6V7AoATb3HPT
H1bROPfoD9Tw6hYASsbwpzGc5sL9X